library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity State_EX_MEM is
    port (
        clk             : in std_logic;
        rst             : in std_logic;
        hazard          : in std_logic;

        
    );
end entity State_EX_MEM;

architecture rtl of State_EX_MEM is
    
begin
    
    
    
end architecture rtl;